PACKAGE FCV IS
    TYPE coloresLED IS (rojo, verde, amarillo, azul, morado, blanco);
	 TYPE posicionesServo IS (abierto, cerrado);
	 TYPE int_array IS array(0 to 5) OF integer;
END PACKAGE;
